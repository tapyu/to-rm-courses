library verilog;
use verilog.vl_types.all;
entity multiplexador2x1_4bits_vlg_vec_tst is
end multiplexador2x1_4bits_vlg_vec_tst;
