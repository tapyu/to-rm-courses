library verilog;
use verilog.vl_types.all;
entity pratica1_vlg_sample_tst is
    port(
        c               : in     vl_logic;
        h               : in     vl_logic;
        p               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end pratica1_vlg_sample_tst;
