library verilog;
use verilog.vl_types.all;
entity pratica1_vlg_check_tst is
    port(
        f               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end pratica1_vlg_check_tst;
