library verilog;
use verilog.vl_types.all;
entity registrador_vlg_vec_tst is
end registrador_vlg_vec_tst;
