library verilog;
use verilog.vl_types.all;
entity pratica1_vlg_vec_tst is
end pratica1_vlg_vec_tst;
