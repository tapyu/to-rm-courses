library verilog;
use verilog.vl_types.all;
entity pratica1 is
    port(
        p               : in     vl_logic;
        c               : in     vl_logic;
        h               : in     vl_logic;
        f               : out    vl_logic
    );
end pratica1;
